*-- interposer PDN spice model 'interposer1' for AC analysis
*-- Total unit cell #: 81 (9x9)

.param cellno=81
.param r_int_cell='1e-3'
.param l_int_cell='1e-10'
.param c_int_cell='1e-11'

xdint_0_0 ndint_x_0_0 ndint_x_1000_0 ndint_y_0_0 ndint_y_0_1000 ndint_xy_0_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_1 ndint_x_1000_0 ndint_x_2000_0 ndint_y_1000_0 ndint_y_1000_1000 ndint_xy_1000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_2 ndint_x_2000_0 ndint_x_3000_0 ndint_y_2000_0 ndint_y_2000_1000 ndint_xy_2000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_3 ndint_x_3000_0 ndint_x_4000_0 ndint_y_3000_0 ndint_y_3000_1000 ndint_xy_3000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_4 ndint_x_4000_0 ndint_x_5000_0 ndint_y_4000_0 ndint_y_4000_1000 ndint_xy_4000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_5 ndint_x_5000_0 ndint_x_6000_0 ndint_y_5000_0 ndint_y_5000_1000 ndint_xy_5000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_6 ndint_x_6000_0 ndint_x_7000_0 ndint_y_6000_0 ndint_y_6000_1000 ndint_xy_6000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_7 ndint_x_7000_0 ndint_x_8000_0 ndint_y_7000_0 ndint_y_7000_1000 ndint_xy_7000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_8 ndint_x_8000_0 ndint_x_9000_0 ndint_y_8000_0 ndint_y_8000_1000 ndint_xy_8000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_0 ndint_x_0_1000 ndint_x_1000_1000 ndint_y_0_1000 ndint_y_0_2000 ndint_xy_0_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_1 ndint_x_1000_1000 ndint_x_2000_1000 ndint_y_1000_1000 ndint_y_1000_2000 ndint_xy_1000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_2 ndint_x_2000_1000 ndint_x_3000_1000 ndint_y_2000_1000 ndint_y_2000_2000 ndint_xy_2000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_3 ndint_x_3000_1000 ndint_x_4000_1000 ndint_y_3000_1000 ndint_y_3000_2000 ndint_xy_3000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_4 ndint_x_4000_1000 ndint_x_5000_1000 ndint_y_4000_1000 ndint_y_4000_2000 ndint_xy_4000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_5 ndint_x_5000_1000 ndint_x_6000_1000 ndint_y_5000_1000 ndint_y_5000_2000 ndint_xy_5000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_6 ndint_x_6000_1000 ndint_x_7000_1000 ndint_y_6000_1000 ndint_y_6000_2000 ndint_xy_6000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_7 ndint_x_7000_1000 ndint_x_8000_1000 ndint_y_7000_1000 ndint_y_7000_2000 ndint_xy_7000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_8 ndint_x_8000_1000 ndint_x_9000_1000 ndint_y_8000_1000 ndint_y_8000_2000 ndint_xy_8000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_0 ndint_x_0_2000 ndint_x_1000_2000 ndint_y_0_2000 ndint_y_0_3000 ndint_xy_0_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_1 ndint_x_1000_2000 ndint_x_2000_2000 ndint_y_1000_2000 ndint_y_1000_3000 ndint_xy_1000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_2 ndint_x_2000_2000 ndint_x_3000_2000 ndint_y_2000_2000 ndint_y_2000_3000 ndint_xy_2000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_3 ndint_x_3000_2000 ndint_x_4000_2000 ndint_y_3000_2000 ndint_y_3000_3000 ndint_xy_3000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_4 ndint_x_4000_2000 ndint_x_5000_2000 ndint_y_4000_2000 ndint_y_4000_3000 ndint_xy_4000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_5 ndint_x_5000_2000 ndint_x_6000_2000 ndint_y_5000_2000 ndint_y_5000_3000 ndint_xy_5000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_6 ndint_x_6000_2000 ndint_x_7000_2000 ndint_y_6000_2000 ndint_y_6000_3000 ndint_xy_6000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_7 ndint_x_7000_2000 ndint_x_8000_2000 ndint_y_7000_2000 ndint_y_7000_3000 ndint_xy_7000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_8 ndint_x_8000_2000 ndint_x_9000_2000 ndint_y_8000_2000 ndint_y_8000_3000 ndint_xy_8000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_0 ndint_x_0_3000 ndint_x_1000_3000 ndint_y_0_3000 ndint_y_0_4000 ndint_xy_0_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_1 ndint_x_1000_3000 ndint_x_2000_3000 ndint_y_1000_3000 ndint_y_1000_4000 ndint_xy_1000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_2 ndint_x_2000_3000 ndint_x_3000_3000 ndint_y_2000_3000 ndint_y_2000_4000 ndint_xy_2000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_3 ndint_x_3000_3000 ndint_x_4000_3000 ndint_y_3000_3000 ndint_y_3000_4000 ndint_xy_3000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_4 ndint_x_4000_3000 ndint_x_5000_3000 ndint_y_4000_3000 ndint_y_4000_4000 ndint_xy_4000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_5 ndint_x_5000_3000 ndint_x_6000_3000 ndint_y_5000_3000 ndint_y_5000_4000 ndint_xy_5000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_6 ndint_x_6000_3000 ndint_x_7000_3000 ndint_y_6000_3000 ndint_y_6000_4000 ndint_xy_6000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_7 ndint_x_7000_3000 ndint_x_8000_3000 ndint_y_7000_3000 ndint_y_7000_4000 ndint_xy_7000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_8 ndint_x_8000_3000 ndint_x_9000_3000 ndint_y_8000_3000 ndint_y_8000_4000 ndint_xy_8000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_0 ndint_x_0_4000 ndint_x_1000_4000 ndint_y_0_4000 ndint_y_0_5000 ndint_xy_0_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_1 ndint_x_1000_4000 ndint_x_2000_4000 ndint_y_1000_4000 ndint_y_1000_5000 ndint_xy_1000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_2 ndint_x_2000_4000 ndint_x_3000_4000 ndint_y_2000_4000 ndint_y_2000_5000 ndint_xy_2000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_3 ndint_x_3000_4000 ndint_x_4000_4000 ndint_y_3000_4000 ndint_y_3000_5000 ndint_xy_3000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_4 ndint_x_4000_4000 ndint_x_5000_4000 ndint_y_4000_4000 ndint_y_4000_5000 ndint_xy_4000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_5 ndint_x_5000_4000 ndint_x_6000_4000 ndint_y_5000_4000 ndint_y_5000_5000 ndint_xy_5000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_6 ndint_x_6000_4000 ndint_x_7000_4000 ndint_y_6000_4000 ndint_y_6000_5000 ndint_xy_6000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_7 ndint_x_7000_4000 ndint_x_8000_4000 ndint_y_7000_4000 ndint_y_7000_5000 ndint_xy_7000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_8 ndint_x_8000_4000 ndint_x_9000_4000 ndint_y_8000_4000 ndint_y_8000_5000 ndint_xy_8000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_0 ndint_x_0_5000 ndint_x_1000_5000 ndint_y_0_5000 ndint_y_0_6000 ndint_xy_0_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_1 ndint_x_1000_5000 ndint_x_2000_5000 ndint_y_1000_5000 ndint_y_1000_6000 ndint_xy_1000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_2 ndint_x_2000_5000 ndint_x_3000_5000 ndint_y_2000_5000 ndint_y_2000_6000 ndint_xy_2000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_3 ndint_x_3000_5000 ndint_x_4000_5000 ndint_y_3000_5000 ndint_y_3000_6000 ndint_xy_3000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_4 ndint_x_4000_5000 ndint_x_5000_5000 ndint_y_4000_5000 ndint_y_4000_6000 ndint_xy_4000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_5 ndint_x_5000_5000 ndint_x_6000_5000 ndint_y_5000_5000 ndint_y_5000_6000 ndint_xy_5000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_6 ndint_x_6000_5000 ndint_x_7000_5000 ndint_y_6000_5000 ndint_y_6000_6000 ndint_xy_6000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_7 ndint_x_7000_5000 ndint_x_8000_5000 ndint_y_7000_5000 ndint_y_7000_6000 ndint_xy_7000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_8 ndint_x_8000_5000 ndint_x_9000_5000 ndint_y_8000_5000 ndint_y_8000_6000 ndint_xy_8000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_0 ndint_x_0_6000 ndint_x_1000_6000 ndint_y_0_6000 ndint_y_0_7000 ndint_xy_0_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_1 ndint_x_1000_6000 ndint_x_2000_6000 ndint_y_1000_6000 ndint_y_1000_7000 ndint_xy_1000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_2 ndint_x_2000_6000 ndint_x_3000_6000 ndint_y_2000_6000 ndint_y_2000_7000 ndint_xy_2000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_3 ndint_x_3000_6000 ndint_x_4000_6000 ndint_y_3000_6000 ndint_y_3000_7000 ndint_xy_3000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_4 ndint_x_4000_6000 ndint_x_5000_6000 ndint_y_4000_6000 ndint_y_4000_7000 ndint_xy_4000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_5 ndint_x_5000_6000 ndint_x_6000_6000 ndint_y_5000_6000 ndint_y_5000_7000 ndint_xy_5000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_6 ndint_x_6000_6000 ndint_x_7000_6000 ndint_y_6000_6000 ndint_y_6000_7000 ndint_xy_6000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_7 ndint_x_7000_6000 ndint_x_8000_6000 ndint_y_7000_6000 ndint_y_7000_7000 ndint_xy_7000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_8 ndint_x_8000_6000 ndint_x_9000_6000 ndint_y_8000_6000 ndint_y_8000_7000 ndint_xy_8000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_0 ndint_x_0_7000 ndint_x_1000_7000 ndint_y_0_7000 ndint_y_0_8000 ndint_xy_0_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_1 ndint_x_1000_7000 ndint_x_2000_7000 ndint_y_1000_7000 ndint_y_1000_8000 ndint_xy_1000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_2 ndint_x_2000_7000 ndint_x_3000_7000 ndint_y_2000_7000 ndint_y_2000_8000 ndint_xy_2000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_3 ndint_x_3000_7000 ndint_x_4000_7000 ndint_y_3000_7000 ndint_y_3000_8000 ndint_xy_3000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_4 ndint_x_4000_7000 ndint_x_5000_7000 ndint_y_4000_7000 ndint_y_4000_8000 ndint_xy_4000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_5 ndint_x_5000_7000 ndint_x_6000_7000 ndint_y_5000_7000 ndint_y_5000_8000 ndint_xy_5000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_6 ndint_x_6000_7000 ndint_x_7000_7000 ndint_y_6000_7000 ndint_y_6000_8000 ndint_xy_6000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_7 ndint_x_7000_7000 ndint_x_8000_7000 ndint_y_7000_7000 ndint_y_7000_8000 ndint_xy_7000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_8 ndint_x_8000_7000 ndint_x_9000_7000 ndint_y_8000_7000 ndint_y_8000_8000 ndint_xy_8000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_0 ndint_x_0_8000 ndint_x_1000_8000 ndint_y_0_8000 ndint_y_0_9000 ndint_xy_0_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_1 ndint_x_1000_8000 ndint_x_2000_8000 ndint_y_1000_8000 ndint_y_1000_9000 ndint_xy_1000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_2 ndint_x_2000_8000 ndint_x_3000_8000 ndint_y_2000_8000 ndint_y_2000_9000 ndint_xy_2000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_3 ndint_x_3000_8000 ndint_x_4000_8000 ndint_y_3000_8000 ndint_y_3000_9000 ndint_xy_3000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_4 ndint_x_4000_8000 ndint_x_5000_8000 ndint_y_4000_8000 ndint_y_4000_9000 ndint_xy_4000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_5 ndint_x_5000_8000 ndint_x_6000_8000 ndint_y_5000_8000 ndint_y_5000_9000 ndint_xy_5000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_6 ndint_x_6000_8000 ndint_x_7000_8000 ndint_y_6000_8000 ndint_y_6000_9000 ndint_xy_6000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_7 ndint_x_7000_8000 ndint_x_8000_8000 ndint_y_7000_8000 ndint_y_7000_9000 ndint_xy_7000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_8 ndint_x_8000_8000 ndint_x_9000_8000 ndint_y_8000_8000 ndint_y_8000_9000 ndint_xy_8000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'


.include 'unitcell.subckt'

rd_ubump2via_0_1 nd_chiplet1_pad_0_1 ndint_y_4000_4000 0.001
rd_ubump2via_0_3 nd_chiplet1_pad_0_3 ndint_y_4000_5000 0.001
rd_ubump2via_0_5 nd_chiplet1_pad_0_5 ndint_y_4000_5000 0.001
rd_ubump2via_0_7 nd_chiplet1_pad_0_7 ndint_y_4000_6000 0.001
rd_ubump2via_0_9 nd_chiplet1_pad_0_9 ndint_y_4000_6000 0.001
rd_ubump2via_1_0 nd_chiplet1_pad_1_0 ndint_y_4000_4000 0.001
rd_ubump2via_1_2 nd_chiplet1_pad_1_2 ndint_y_4000_4000 0.001
rd_ubump2via_1_4 nd_chiplet1_pad_1_4 ndint_y_4000_5000 0.001
rd_ubump2via_1_6 nd_chiplet1_pad_1_6 ndint_y_4000_5000 0.001
rd_ubump2via_1_8 nd_chiplet1_pad_1_8 ndint_y_4000_6000 0.001
rd_ubump2via_2_1 nd_chiplet1_pad_2_1 ndint_y_4000_4000 0.001
rd_ubump2via_2_3 nd_chiplet1_pad_2_3 ndint_y_4000_5000 0.001
rd_ubump2via_2_5 nd_chiplet1_pad_2_5 ndint_y_4000_5000 0.001
rd_ubump2via_2_7 nd_chiplet1_pad_2_7 ndint_y_4000_6000 0.001
rd_ubump2via_2_9 nd_chiplet1_pad_2_9 ndint_y_4000_6000 0.001
rd_ubump2via_3_0 nd_chiplet1_pad_3_0 ndint_y_5000_4000 0.001
rd_ubump2via_3_2 nd_chiplet1_pad_3_2 ndint_y_5000_4000 0.001
rd_ubump2via_3_4 nd_chiplet1_pad_3_4 ndint_y_5000_5000 0.001
rd_ubump2via_3_6 nd_chiplet1_pad_3_6 ndint_y_5000_5000 0.001
rd_ubump2via_3_8 nd_chiplet1_pad_3_8 ndint_y_5000_6000 0.001
rd_ubump2via_4_1 nd_chiplet1_pad_4_1 ndint_y_5000_4000 0.001
rd_ubump2via_4_3 nd_chiplet1_pad_4_3 ndint_y_5000_5000 0.001
rd_ubump2via_4_5 nd_chiplet1_pad_4_5 ndint_y_5000_5000 0.001
rd_ubump2via_4_7 nd_chiplet1_pad_4_7 ndint_y_5000_6000 0.001
rd_ubump2via_4_9 nd_chiplet1_pad_4_9 ndint_y_5000_6000 0.001
rd_ubump2via_5_0 nd_chiplet1_pad_5_0 ndint_y_5000_4000 0.001
rd_ubump2via_5_2 nd_chiplet1_pad_5_2 ndint_y_5000_4000 0.001
rd_ubump2via_5_4 nd_chiplet1_pad_5_4 ndint_y_5000_5000 0.001
rd_ubump2via_5_6 nd_chiplet1_pad_5_6 ndint_y_5000_5000 0.001
rd_ubump2via_5_8 nd_chiplet1_pad_5_8 ndint_y_5000_6000 0.001
rd_ubump2via_6_1 nd_chiplet1_pad_6_1 ndint_y_5000_4000 0.001
rd_ubump2via_6_3 nd_chiplet1_pad_6_3 ndint_y_5000_5000 0.001
rd_ubump2via_6_5 nd_chiplet1_pad_6_5 ndint_y_5000_5000 0.001
rd_ubump2via_6_7 nd_chiplet1_pad_6_7 ndint_y_5000_6000 0.001
rd_ubump2via_6_9 nd_chiplet1_pad_6_9 ndint_y_5000_6000 0.001
rd_ubump2via_7_0 nd_chiplet1_pad_7_0 ndint_y_6000_4000 0.001
rd_ubump2via_7_2 nd_chiplet1_pad_7_2 ndint_y_6000_4000 0.001
rd_ubump2via_7_4 nd_chiplet1_pad_7_4 ndint_y_6000_5000 0.001
rd_ubump2via_7_6 nd_chiplet1_pad_7_6 ndint_y_6000_5000 0.001
rd_ubump2via_7_8 nd_chiplet1_pad_7_8 ndint_y_6000_6000 0.001
rd_ubump2via_8_1 nd_chiplet1_pad_8_1 ndint_y_6000_4000 0.001
rd_ubump2via_8_3 nd_chiplet1_pad_8_3 ndint_y_6000_5000 0.001
rd_ubump2via_8_5 nd_chiplet1_pad_8_5 ndint_y_6000_5000 0.001
rd_ubump2via_8_7 nd_chiplet1_pad_8_7 ndint_y_6000_6000 0.001
rd_ubump2via_8_9 nd_chiplet1_pad_8_9 ndint_y_6000_6000 0.001
rd_ubump2via_9_0 nd_chiplet1_pad_9_0 ndint_y_6000_4000 0.001
rd_ubump2via_9_2 nd_chiplet1_pad_9_2 ndint_y_6000_4000 0.001
rd_ubump2via_9_4 nd_chiplet1_pad_9_4 ndint_y_6000_5000 0.001
rd_ubump2via_9_6 nd_chiplet1_pad_9_6 ndint_y_6000_5000 0.001
rd_ubump2via_9_8 nd_chiplet1_pad_9_8 ndint_y_6000_6000 0.001

*-- chiplet instance [0]: chiplet1
xchiplet_chiplet1
+nd_chiplet1_pad_0_1
+nd_chiplet1_pad_0_3
+nd_chiplet1_pad_0_5
+nd_chiplet1_pad_0_7
+nd_chiplet1_pad_0_9
+nd_chiplet1_pad_1_0
+nd_chiplet1_pad_1_2
+nd_chiplet1_pad_1_4
+nd_chiplet1_pad_1_6
+nd_chiplet1_pad_1_8
+nd_chiplet1_pad_2_1
+nd_chiplet1_pad_2_3
+nd_chiplet1_pad_2_5
+nd_chiplet1_pad_2_7
+nd_chiplet1_pad_2_9
+nd_chiplet1_pad_3_0
+nd_chiplet1_pad_3_2
+nd_chiplet1_pad_3_4
+nd_chiplet1_pad_3_6
+nd_chiplet1_pad_3_8
+nd_chiplet1_pad_4_1
+nd_chiplet1_pad_4_3
+nd_chiplet1_pad_4_5
+nd_chiplet1_pad_4_7
+nd_chiplet1_pad_4_9
+nd_chiplet1_pad_5_0
+nd_chiplet1_pad_5_2
+nd_chiplet1_pad_5_4
+nd_chiplet1_pad_5_6
+nd_chiplet1_pad_5_8
+nd_chiplet1_pad_6_1
+nd_chiplet1_pad_6_3
+nd_chiplet1_pad_6_5
+nd_chiplet1_pad_6_7
+nd_chiplet1_pad_6_9
+nd_chiplet1_pad_7_0
+nd_chiplet1_pad_7_2
+nd_chiplet1_pad_7_4
+nd_chiplet1_pad_7_6
+nd_chiplet1_pad_7_8
+nd_chiplet1_pad_8_1
+nd_chiplet1_pad_8_3
+nd_chiplet1_pad_8_5
+nd_chiplet1_pad_8_7
+nd_chiplet1_pad_8_9
+nd_chiplet1_pad_9_0
+nd_chiplet1_pad_9_2
+nd_chiplet1_pad_9_4
+nd_chiplet1_pad_9_6
+nd_chiplet1_pad_9_8
+chiplet1
.include 'chiplet1_tr_new.subckt'

*-- tsv array
xdint_tsv_0_1 ndint_tsv_0_1 ndint_bump_0_1 int_tsv
xdint_tsv_0_3 ndint_tsv_0_3 ndint_bump_0_3 int_tsv
xdint_tsv_1_0 ndint_tsv_1_0 ndint_bump_1_0 int_tsv
xdint_tsv_1_2 ndint_tsv_1_2 ndint_bump_1_2 int_tsv
xdint_tsv_1_4 ndint_tsv_1_4 ndint_bump_1_4 int_tsv
xdint_tsv_2_1 ndint_tsv_2_1 ndint_bump_2_1 int_tsv
xdint_tsv_2_3 ndint_tsv_2_3 ndint_bump_2_3 int_tsv
xdint_tsv_3_0 ndint_tsv_3_0 ndint_bump_3_0 int_tsv
xdint_tsv_3_2 ndint_tsv_3_2 ndint_bump_3_2 int_tsv
xdint_tsv_3_4 ndint_tsv_3_4 ndint_bump_3_4 int_tsv
xdint_tsv_4_1 ndint_tsv_4_1 ndint_bump_4_1 int_tsv
xdint_tsv_4_3 ndint_tsv_4_3 ndint_bump_4_3 int_tsv
.include 'int_tsv.subckt'

*-- tsv to via
rdint_tsv2via_0_1 ndint_tsv_0_1 ndint_y_2000_3000 0.001
rdint_tsv2via_0_3 ndint_tsv_0_3 ndint_xy_2000_7000 0.001
rdint_tsv2via_1_0 ndint_tsv_1_0 ndint_y_3000_2000 0.001
rdint_tsv2via_1_2 ndint_tsv_1_2 ndint_y_3000_5000 0.001
rdint_tsv2via_1_4 ndint_tsv_1_4 ndint_xy_3000_8000 0.001
rdint_tsv2via_2_1 ndint_tsv_2_1 ndint_y_5000_3000 0.001
rdint_tsv2via_2_3 ndint_tsv_2_3 ndint_y_5000_7000 0.001
rdint_tsv2via_3_0 ndint_tsv_3_0 ndint_xy_7000_2000 0.001
rdint_tsv2via_3_2 ndint_tsv_3_2 ndint_y_7000_5000 0.001
rdint_tsv2via_3_4 ndint_tsv_3_4 ndint_y_7000_8000 0.001
rdint_tsv2via_4_1 ndint_tsv_4_1 ndint_xy_8000_3000 0.001
rdint_tsv2via_4_3 ndint_tsv_4_3 ndint_y_8000_7000 0.001

*-- tsv bump array to pkg
rdint_tsv_0_1 ndint_bump_0_1 nd_pkg_pad 0.001
rdint_tsv_0_3 ndint_bump_0_3 nd_pkg_pad 0.001
rdint_tsv_1_0 ndint_bump_1_0 nd_pkg_pad 0.001
rdint_tsv_1_2 ndint_bump_1_2 nd_pkg_pad 0.001
rdint_tsv_1_4 ndint_bump_1_4 nd_pkg_pad 0.001
rdint_tsv_2_1 ndint_bump_2_1 nd_pkg_pad 0.001
rdint_tsv_2_3 ndint_bump_2_3 nd_pkg_pad 0.001
rdint_tsv_3_0 ndint_bump_3_0 nd_pkg_pad 0.001
rdint_tsv_3_2 ndint_bump_3_2 nd_pkg_pad 0.001
rdint_tsv_3_4 ndint_bump_3_4 nd_pkg_pad 0.001
rdint_tsv_4_1 ndint_bump_4_1 nd_pkg_pad 0.001
rdint_tsv_4_3 ndint_bump_4_3 nd_pkg_pad 0.001

*-- pkg instances
xpkg_vdd vdd_pkg nd_pkg_pad pkg_model
.include 'pkg.subckt'

*-- pcb instances
xpcb_vdd vdd vdd_pkg pcb_model
.include 'pcb.subckt'
*--.include 'vdd_decap.1'

*-- external power source
vdd vdd 0 1
.tran 1.000000e-11 1.000000e-08
.end
